-- Biên dịch chương trình và testbench:
--   ghdl -a InstructionMemory.vhd
--   ghdl -a InstructionMemory_tb.vhd
--
-- Chạy mô phỏng:
--   ghdl -e InstructionMemory_tb
--   ghdl -r InstructionMemory_tb --vcd=imem_wave.vcd
--   gtkwave imem_wave.vcd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;   

entity InstructionMemory is
    port(
        Address     : in  STD_LOGIC_VECTOR(31 downto 0); -- Địa chỉ byte từ PC
        Instruction : out STD_LOGIC_VECTOR(31 downto 0)  -- Lệnh 32 bit
    );
end entity;

architecture Behavioral of InstructionMemory is

    -----------------------------------------------------------
    -- ROM: Mảng hằng các lệnh MIPS (32-bit)
    -----------------------------------------------------------
    type ROM_ARRAY is array (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
    -- Vị trí nhập lệnh vào ROM
    constant ROM : ROM_ARRAY := (
        -- 0: addi $t0, $zero, 10      ($t0 = 10)
        0 => x"2008000A", 
        
        -- 1: j 4                      (Nhảy đến index 4)
        -- Opcode j=000010. Target=4. Hex: 08000004
        1 => x"08000004", 
        
        -- 2: addi $t0, $zero, 99      (TRAP: Nếu j sai, $t0 = 99)
        2 => x"20080063",
        
        -- 3: addi $t0, $zero, 99      (TRAP: Lệnh rác)
        3 => x"20080063", 
        
        -- 4: Label_Target_J: addi $t1, $zero, 20  ($t1 = 20)
        4 => x"20090014",
        
        -- 5: jal 8                    (Nhảy đến index 8, lưu PC+4 vào $31)
        -- Opcode jal=000011. Target=8. Hex: 0C000008
        -- PC hiện tại là 5*4=20. PC+4 = 24 (0x18). Vậy $31 sẽ bằng 24.
        5 => x"0C000008",
        
        -- 6: addi $t2, $zero, 99      (TRAP: Nếu jal sai, $t2 = 99)
        6 => x"200A0063",
        
        -- 7: addi $t2, $zero, 99      (TRAP: Lệnh rác)
        7 => x"200A0063",
        
        -- 8: Label_Target_JAL: addi $t3, $ra, 0   ($t3 = $ra)
        -- Để kiểm tra xem $ra có đúng là 24 (0x18) không.
        8 => x"23EB0000",
        
        -- 9: j 9                      (Vòng lặp vô tận để dừng chương trình)
        9 => x"08000009",
        others => x"00000000"
    );

begin

    -----------------------------------------------------------
    -- Xuất lệnh tương ứng với Address(31 downto 2) 
    -- Bỏ 2 bít cuối vì 2 bít cuối là chỉ tới vị trí thứ mấy trong từ 4 byte
    -- Quy trình: hex => nhị phân => lấy 31 đến 2 => chuyển sang số nguyên 
    -- Thực hiện dịch phải 2 bit (tương ứng với việc nhân 4 byte) để chuyển địa chỉ byte thành chỉ số word trong ROM
    -----------------------------------------------------------
    Instruction <= ROM(to_integer(unsigned(Address(31 downto 2))));

end architecture;
