-- Biên dịch chương trình và testbench:
--   ghdl -a InstructionMemory.vhd
--   ghdl -a InstructionMemory_tb.vhd
--
-- Chạy mô phỏng:
--   ghdl -e InstructionMemory_tb
--   ghdl -r InstructionMemory_tb --vcd=imem_wave.vcd
--   gtkwave imem_wave.vcd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;   

entity InstructionMemory is
    port(
        Address     : in  STD_LOGIC_VECTOR(31 downto 0); -- Địa chỉ byte từ PC
        Instruction : out STD_LOGIC_VECTOR(31 downto 0)  -- Lệnh 32 bit
    );
end entity;

architecture Behavioral of InstructionMemory is

    -----------------------------------------------------------
    -- ROM: Mảng hằng các lệnh MIPS (32-bit)
    -----------------------------------------------------------
    type ROM_ARRAY is array (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
    -- Vị trí nhập lệnh vào ROM
    constant ROM : ROM_ARRAY := (
        -- Test beq và bne
        0 => x"20080005",  -- addi $t0, $zero, 5     # $t0 = 5
        1 => x"20090005",  -- addi $t1, $zero, 5     # $t1 = 5
        2 => x"200A0003",  -- addi $t2, $zero, 3     # $t2 = 3
        3 => x"11090002",  -- beq $t0, $t1, label1   # branch nếu $t0 == $t1 (sẽ nhảy)
        4 => x"200B0001",  -- addi $t3, $zero, 1     # $t3 = 1 (bị bỏ qua)
        5 => x"200B0002",  -- addi $t3, $zero, 2     # $t3 = 2 (bị bỏ qua)
        6 => x"200C00FF",  -- label1: addi $t4, $zero, 255  # $t4 = 255
        7 => x"150A0002",  -- bne $t0, $t2, label2   # branch nếu $t0 != $t2 (sẽ nhảy)
        8 => x"200D0001",  -- addi $t5, $zero, 1     # $t5 = 1 (bị bỏ qua)
        9 => x"200D0002",  -- addi $t5, $zero, 2     # $t5 = 2 (bị bỏ qua)
        10 => x"200E00AA", -- label2: addi $t6, $zero, 170  # $t6 = 170
        others => x"00000000"
    );

begin

    -----------------------------------------------------------
    -- Xuất lệnh tương ứng với Address(31 downto 2) 
    -- Bỏ 2 bít cuối vì 2 bít cuối là chỉ tới vị trí thứ mấy trong từ 4 byte
    -- Quy trình: hex => nhị phân => lấy 31 đến 2 => chuyển sang số nguyên 
    -- Thực hiện dịch phải 2 bit (tương ứng với việc nhân 4 byte) để chuyển địa chỉ byte thành chỉ số word trong ROM
    -----------------------------------------------------------
    Instruction <= ROM(to_integer(unsigned(Address(31 downto 2))));

end architecture;
