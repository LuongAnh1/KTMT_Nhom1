-- B1: Nhập lệnh dưới dạng mã hex vào Instruction Memory (ROM)
-- B2: Kết nối các khối để tạo thành CPU đơn chu kỳ hoàn chỉnh
-- Biên dịch CPU đơn chu kỳ (Nạp dữ liệu vào thanh ghi và bắt đầu chạy ở giây thứu 300ns):
-- ghdl -a BrentKung_16.vhd BrentKung_32.vhd
-- ghdl -a PC.vhd InstructionMemory.vhd CU.vhd RegisterFile.vhd ALUControl.vhd ALU.vhd DataMemory.vhd MUX_WriteBack.vhd CPU.vhd CPU_tb.vhd
-- ghdl -e SingleCycleCPU_tb
-- ghdl -r SingleCycleCPU_tb --vcd=singlecpu.vcd --stop-time=300ns
-- gtkwave singlecpu.vcd

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SingleCycleCPU IS
    PORT (
        clk, reset : IN STD_LOGIC;

        -- Phần hỗ trợ test bench
        -- Tín hiệu để ghi dữ liệu cho thanh ghi từ test bench
        dbg_write_enable : in std_logic := '0'; 
        -- '1' thì test bench được ghi, '0' thì CPU bình thường ghi
        dbg_write_reg    : in std_logic_vector(4 downto 0) := (others => '0'); 
        -- Địa chỉ thanh ghi muốn ghi 
        dbg_write_data   : in std_logic_vector(31 downto 0) := (others => '0');
        -- Dữ liệu mà testbench muốn nạp vào thanh ghi
        dbg_read_reg     : in std_logic_vector(4 downto 0) := (others => '0');
        -- Testbench yêu cầu đọc nội dung của thanh ghi nào
        dbg_read_data    : out std_logic_vector(31 downto 0) 
        -- Xuất giá trị thanh ghi ra test bench, không ảnh hưởng đến hoạt động CPU
    );
END ENTITY;

ARCHITECTURE behavior OF SingleCycleCPU IS

    -- ==== Tín hiệu liên kết các khối ====
    SIGNAL PC_in, PC_out             : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL Instruction               : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL ReadData1, ReadData2      : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL SignImm                   : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL ALUResult, MemReadData    : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL WriteDataReg              : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL Zero                      : STD_LOGIC;
    SIGNAL ALUControlSig             : STD_LOGIC_VECTOR(3 DOWNTO 0);

    -- Tín hiệu cho các MUX
    SIGNAL WriteRegAddr              : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL ALU_B                     : STD_LOGIC_VECTOR(31 DOWNTO 0);

    -- Control Unit outputs
    SIGNAL RegDst, ALUSrc, MemToReg, RegWrite, MemRead, MemWrite, Branch : STD_LOGIC;
    SIGNAL ALUOp                     : STD_LOGIC_VECTOR(1 DOWNTO 0);

    signal RF_WriteReg  : std_logic_vector(4 downto 0);
    signal RF_WriteData : std_logic_vector(31 downto 0);
    signal RF_RegWrite  : std_logic;

BEGIN
    
    ------------------------------------------------------------------------
    -- 1. Program Counter
    ------------------------------------------------------------------------
    PC_inst: ENTITY work.PC
        PORT MAP (
            clk => clk, -- xung nhịp cho PC (in)
            reset => reset, -- tín hiệu reset cho PC (in)
            PC_in => PC_in, -- địa chỉ lệnh tiếp theo (in)
            PC_out => PC_out -- địa chỉ lệnh hiện tại (out)
        );

    ------------------------------------------------------------------------
    -- 2. Instruction Memory
    ------------------------------------------------------------------------
    IM_inst: ENTITY work.InstructionMemory
        PORT MAP (
            Address => PC_out, -- địa chỉ lệnh từ PC (in)
            Instruction => Instruction -- lệnh ra (out)
        );

    ------------------------------------------------------------------------
    -- 3. Control Unit
    ------------------------------------------------------------------------
    CU_inst: ENTITY work.ControlUnit
        PORT MAP (
            opcode    => Instruction(31 DOWNTO 26),
            RegDst    => RegDst, -- tín hiệu chọn WriteReg
            ALUSrc    => ALUSrc, -- tín hiệu chọn ALU input B (ReadData2 hoặc SignImm)
            MemToReg  => MemToReg, -- tín hiệu chọn dữ liệu ghi vào Register File (ALUResult hoặc MemReadData)
            RegWrite  => RegWrite, -- tín hiệu cho phép ghi vào Register File
            MemRead   => MemRead, -- tín hiệu đọc từ Data Memory
            MemWrite  => MemWrite, -- tín hiệu ghi vào Data Memory
            Branch    => Branch, -- tín hiệu nhánh
            ALUOp     => ALUOp -- tín hiệu điều khiển ALU
        );


    ------------------------------------------------------------------------
    -- Sign Extend (16-bit immediate -> 32-bit)
    ------------------------------------------------------------------------
    SignImm <= (31 DOWNTO 16 => Instruction(15)) & Instruction(15 DOWNTO 0);

    ------------------------------------------------------------------------
    -- MUX RegDst (chọn WriteReg: rd hoặc rt)
    ------------------------------------------------------------------------
    -- Nếu RegDst = 1 ~ R-type thì chọn rd (Instruction[15:11])
    -- Ngược lại chọn rt ~ I-type (Instruction[20:16])
    WriteRegAddr <= Instruction(15 DOWNTO 11) WHEN RegDst = '1' 
                    ELSE Instruction(20 DOWNTO 16);


    ------------------------------------------------------------------------
    -- 4. Register File
    ------------------------------------------------------------------------
    -- Nếu debug đang bật => test bench điều khiển ghi thanh ghi (register file)
    -- Ngược lại CPU hoạt động bình thường

    RF_RegWrite  <= dbg_write_enable or RegWrite;
    -- Nếu testbench bật debug (dbg_write_enable = 1) → Register File sẽ cho phép ghi
    -- Nếu CPU yêu cầu ghi (RegWrite = 1) → Register File ghi theo CPU
    -- Nếu cả hai đều 0 → Register File không ghi

    RF_WriteReg  <= dbg_write_reg  when dbg_write_enable = '1'
                    else WriteRegAddr;
    -- Nếu debug bật:
    --     Testbench chọn thanh ghi cần ghi qua dbg_write_reg
    --     CPU bị vô hiệu hóa, không chọn được
    -- Nếu debug tắt:CPU chọn thanh ghi đích bình thường (WriteRegAddr = rd hoặc rt)

    RF_WriteData <= dbg_write_data when dbg_write_enable = '1'
                    else WriteDataReg;
    -- Debug bật: Testbench nạp giá trị trực tiếp vào thanh ghi (dbg_write_data)
    -- Debug tắt: CPU ghi dữ liệu tính từ MUX WriteBack (WriteDataReg)

    RF_inst: ENTITY work.RegisterFile
        PORT MAP (
            clk        => clk,
            RegWrite   => RF_RegWrite, -- tín hiệu từ Control Unit (Cho phép ghi hay không) (in)
            ReadReg1   => Instruction(25 downto 21),
            ReadReg2   => Instruction(20 downto 16),
            WriteReg   => RF_WriteReg,
            WriteData  => RF_WriteData,
            ReadData1  => ReadData1,
            ReadData2  => ReadData2
            -- clk        => clk, -- xung nhịp cho Register File (in)
            -- RegWrite   => RegWrite, -- tín hiệu từ Control Unit (Cho phép ghi hay không) (in)
            -- ReadReg1   => Instruction(25 DOWNTO 21), -- rs: thanh ghi nguồn 1 (in)
            -- ReadReg2   => Instruction(20 DOWNTO 16), -- rt: thanh ghi nguồn 2 (in)
            -- WriteReg   => WriteRegAddr, -- tín hiệu từ MUX RegDst (chọn rd hoặc rt) (in)
            -- WriteData  => WriteDataReg, -- dữ liệu ghi vào thanh ghi đích (in)
            -- ReadData1  => ReadData1, -- dữ liệu đọc từ thanh ghi nguồn 1 (out)
            -- ReadData2  => ReadData2 -- dữ liệu đọc từ thanh ghi nguồn 2 (out)
        );

    
    ------------------------------------------------------------------------
    -- MUX ALUSrc (chọn ALU input B: ReadData2 ~ rd (R-type) hoặc SignImm ~ immediate (I-type))
    ------------------------------------------------------------------------
    ALU_B <= SignImm WHEN ALUSrc = '1' ELSE ReadData2;


    ------------------------------------------------------------------------
    -- 5. ALU Control
    ------------------------------------------------------------------------
    ALUC_inst: ENTITY work.ALUCO
        PORT MAP (
            ALUOp      => ALUOp, -- tín hiệu từ Control Unit (in)
            funct      => Instruction(5 DOWNTO 0), -- phần funct của lệnh R-type (in)
            ALUControl => ALUControlSig -- tín hiệu điều khiển ALU (out)
        );

    ------------------------------------------------------------------------
    -- 6. ALU
    ------------------------------------------------------------------------
    ALU_inst: ENTITY work.ALU
        PORT MAP (
            A           => ReadData1, -- từ Register File (in)
            B           => ALU_B,   -- từ MUX ALUSrc (ReadData2 hoặc Immediate) (in)
            ALUControl  => ALUControlSig, -- từ ALU Control (in)
            Result      => ALUResult, -- kết quả ALU (out)
            Zero        => Zero -- tín hiệu Zero (out)
        );

    ------------------------------------------------------------------------
    -- 7. Data Memory
    ------------------------------------------------------------------------
    DM_inst: ENTITY work.DataMemory
        PORT MAP (
            clk        => clk, -- xung nhịp cho Data Memory (in)
            MemRead    => MemRead, -- Cho phép đọc từ Data Memory (in)
            MemWrite   => MemWrite, -- Cho phép ghi vào Data Memory (in)
            Address    => ALUResult, -- địa chỉ ô nhớ cần đọc/ghi từ ALU (in)
            WriteData  => ReadData2, -- dữ liệu cần ghi vào Data Memory từ Register File (in)
            ReadData   => MemReadData -- dữ liệu đọc từ Data Memory (out)
        );

    ------------------------------------------------------------------------
    -- 8. MUX WriteBack
    -- Chức năng: Chọn dữ liệu ghi vào Register File (ALUResult hoặc MemReadData)
    ------------------------------------------------------------------------
    WB_mux: ENTITY work.MUX_WriteBack
        PORT MAP (
            ALUResult  => ALUResult, -- kết quả từ ALU (in)
            ReadData   => MemReadData, -- dữ liệu từ Data Memory (in)
            MemToReg   => MemToReg, -- tín hiệu từ Control Unit (in)
            WriteData  => WriteDataReg -- dữ liệu ghi vào Register File (out)
        );

    ------------------------------------------------------------------------
    -- 9. PC Update (tăng +4 đơn giản)
    ------------------------------------------------------------------------
    PC_in <= STD_LOGIC_VECTOR(unsigned(PC_out) + 4);

END ARCHITECTURE;
