                    ┌───────────────────────────────┐
                    │           Control Unit        │
                    │                               │
                    │  ┌───────────────┐            │
                    │  │  ALU Control  │◄───────────┤
                    │  └───────────────┘            │
                    │ RegDst, ALUSrc, MemtoReg,     │
                    │ RegWrite, MemRead, MemWrite,  │
                    │ Branch, PCSrc, ALUOp          │
                    └──────────────┬────────────────┘
                                   │
                                   ▼
 ┌─────────────┐       ┌─────────────────────┐       ┌─────────────┐
 │ Program     │       │ Instruction Memory  │       │  Register   │
 │ Counter (PC)│──►───▶│  (ROM chứa lệnh)   │──►───▶│   File      │
 │             │       │   Instr[31:0]      │        │ (rs, rt, rd)│
 └─────────────┘       └─────────────────────┘       └─────────────┘
       ▲                         │                        │
       │                         │                        │
       │                         ▼                        ▼
       │               ┌────────────────┐       ┌────────────────┐
       │               │ Sign Extend    │       │     MUX        │◄── RegDst
       │               │ (Imm[15:0]→32b)│       └────────────────┘
       │               └────────────────┘               │
       │                         │                     ▼
       │                         └──────┐        ┌────────────┐
       │                                ▼        │    ALU     │
       │                           ┌──────────┐  │            │
       │                           │  MUX     │◄─┤ ALUSrc     │
       │                           └──────────┘  └────────────┘
       │                                │              │
       │                                ▼              ▼
       │                          ┌────────────────────────┐
       │                          │     Data Memory        │
       │                          │  (RAM, LW/SW access)  │
       │                          └────────────────────────┘
       │                                │
       │                                ▼
       │                         ┌─────────────┐
       │                         │     MUX     │◄── MemtoReg
       │                         └─────────────┘
       │                                │
       │                                ▼
       │                         ┌─────────────┐
       │                         │ Write Back  │
       │                         └─────────────┘
       │
       ▼
 ┌──────────────────────┐
 │ PC Update Logic      │
 │ (Adder, Branch, MUX) │
 └──────────────────────┘
             │
             ▼
            PCNext ──► (đưa về PC đầu chu kỳ sau)

-----------------------------------------------------------------------------------------------
-- Module và các tín hiệu điều khiển chính 
-- Sign Extend: Mở rộng immediate từ 16 lên 32 bit
-- Control Unit: Tạo các tín hiệu điều khiển dựa trên opcode và funct
-- Register File: (Điều khiển: RegWrite)
-- ALU: (Điều khiển: ALUSrc)
-- Data Memory: Đọc/Ghi bộ nhớ dữ liệu (Điều khiển: MemRead, MemWrite)
-- Mux: Chọn giữa các nguồn dữ liệu khác nhau (Điều khiển: RegDst, ALUSrc, MemtoReg, PCSrc)
-- Branch Add: Tính địa chỉ tiếp theo hoặc nhánh (Điều khiển: PCSrc)
                ┌────────────────────────────────────────────────┐
                │                     CPU                        │
                └────────────────────────────────────────────────┘
                                ▲
                                │ PCSrc
                                │
                   ┌────────────┴────────────┐
                   │                         │
                   ▼                         │
        ┌───────────────────┐                │
        │Program Counter(PC)│◄─────────────┐ │
        └───────┬───────────┘              │ │
                │ PC + 4                   │ │
                ▼                          │ │
        ┌──────────────────┐               │ │
        │ Instruction Mem  │               │ │
        └───────┬──────────┘               │ │
                │ Instruction[31:0]        │ │
                ▼                          │ │
        ┌──────────────────────────────────────────┐
        │                 Control Unit             │
        ├──────────────────────────────────────────┤
        │ RegDst │ ALUSrc │ MemtoReg │ RegWrite    │
        │ MemRead│ MemWrite│ Branch  │ ALUOp[1:0]  │
        └──────────────────────────────────────────┘
                │
                │ Control Signals
                ▼
        ┌─────────────────────────────┐
        │   Register File             │
        │  ┌───────────────────────┐  │
        │  │ rs ──►│               │  │
        │  │ rt ──►│   Read Ports  │  │
        │  │ rd ◄──│   Write Port  │  │
        │  └───────────────────────┘  │
        └────────┬──────────────┬─────┘
                 │              │
                 ▼              ▼
   ┌─────────────────────┐  ┌───────────────┐
   │Sign-Extend (16->32b)|  │   ALU Control │
   └────────────┬────────┘  └──────┬────────┘
                │                  │
                ▼                  ▼
        ┌──────────────────────────────────────────┐
        │                 ALU                      │
        │   ┌──────────────────────────────────┐   │
        │   │  ALUResult = (A op B)            │   │
        │   └──────────────────────────────────┘   │
        └──────┬──────────────┬────────────────────┘
               │              │
               ▼              ▼
     ┌──────────────────┐   ┌──────────────────┐
     │   Data Memory    │ ->│   Mux (MemtoReg) │
     └──────────────────┘   └──────────────────┘
               │                     │
               │                     ▼
               │              Write Back to Register File
               │
               ▼
          ┌───────────┐
          │   PC + 4  │
          └────┬──────┘
               │
               ▼
        ┌───────────────┐
        │ Branch Add    │
        └────┬──────────┘
             │
             ▼
          Mux (PCSrc) ───► Next PC

-----------------------------------------------------------------------------------------------
